vbhfl
